//Copyright (C)2014-2023 Gowin Semiconductor Corporation.
//All rights reserved.
//File Title: IP file
//Tool Version: V1.9.9 (64-bit)
//Part Number: GW2A-LV18PG256C8/I7
//Device: GW2A-18
//Device Version: C
//Created Time: Sat Sep 27 07:26:32 2025

module blk_mem_gen_4 (douta, doutb, clka, ocea, cea, reseta, wrea, clkb, oceb, ceb, resetb, wreb, ada, dina, adb, dinb);

output [7:0] douta;
output [7:0] doutb;
input clka;
input ocea;
input cea;
input reseta;
input wrea;
input clkb;
input oceb;
input ceb;
input resetb;
input wreb;
input [14:0] ada;
input [7:0] dina;
input [14:0] adb;
input [7:0] dinb;

wire [14:0] dpb_inst_0_douta_w;
wire [0:0] dpb_inst_0_douta;
wire [14:0] dpb_inst_0_doutb_w;
wire [0:0] dpb_inst_0_doutb;
wire [14:0] dpb_inst_1_douta_w;
wire [1:1] dpb_inst_1_douta;
wire [14:0] dpb_inst_1_doutb_w;
wire [1:1] dpb_inst_1_doutb;
wire [14:0] dpb_inst_2_douta_w;
wire [2:2] dpb_inst_2_douta;
wire [14:0] dpb_inst_2_doutb_w;
wire [2:2] dpb_inst_2_doutb;
wire [14:0] dpb_inst_3_douta_w;
wire [3:3] dpb_inst_3_douta;
wire [14:0] dpb_inst_3_doutb_w;
wire [3:3] dpb_inst_3_doutb;
wire [11:0] dpb_inst_4_douta_w;
wire [3:0] dpb_inst_4_douta;
wire [11:0] dpb_inst_4_doutb_w;
wire [3:0] dpb_inst_4_doutb;
wire [14:0] dpb_inst_5_douta_w;
wire [4:4] dpb_inst_5_douta;
wire [14:0] dpb_inst_5_doutb_w;
wire [4:4] dpb_inst_5_doutb;
wire [14:0] dpb_inst_6_douta_w;
wire [5:5] dpb_inst_6_douta;
wire [14:0] dpb_inst_6_doutb_w;
wire [5:5] dpb_inst_6_doutb;
wire [14:0] dpb_inst_7_douta_w;
wire [6:6] dpb_inst_7_douta;
wire [14:0] dpb_inst_7_doutb_w;
wire [6:6] dpb_inst_7_doutb;
wire [14:0] dpb_inst_8_douta_w;
wire [7:7] dpb_inst_8_douta;
wire [14:0] dpb_inst_8_doutb_w;
wire [7:7] dpb_inst_8_doutb;
wire [11:0] dpb_inst_9_douta_w;
wire [7:4] dpb_inst_9_douta;
wire [11:0] dpb_inst_9_doutb_w;
wire [7:4] dpb_inst_9_doutb;
wire dff_q_0;
wire dff_q_1;
wire dff_q_2;
wire cea_w;
wire ceb_w;
wire gw_gnd;

assign cea_w = ~wrea & cea;
assign ceb_w = ~wreb & ceb;
assign gw_gnd = 1'b0;

DPB dpb_inst_0 (
    .DOA({dpb_inst_0_douta_w[14:0],dpb_inst_0_douta[0]}),
    .DOB({dpb_inst_0_doutb_w[14:0],dpb_inst_0_doutb[0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[0]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[0]})
);

defparam dpb_inst_0.READ_MODE0 = 1'b0;
defparam dpb_inst_0.READ_MODE1 = 1'b1;
defparam dpb_inst_0.WRITE_MODE0 = 2'b00;
defparam dpb_inst_0.WRITE_MODE1 = 2'b00;
defparam dpb_inst_0.BIT_WIDTH_0 = 1;
defparam dpb_inst_0.BIT_WIDTH_1 = 1;
defparam dpb_inst_0.BLK_SEL_0 = 3'b000;
defparam dpb_inst_0.BLK_SEL_1 = 3'b000;
defparam dpb_inst_0.RESET_MODE = "SYNC";
defparam dpb_inst_0.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFF053FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFF053FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFF11477FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFF845CF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_06 = 256'h0000FFFFFFFFFFFFFFF0442E2DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_07 = 256'h0000FFFFFFFFFFFFFFFD47150FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_08 = 256'h0000FFFFFFFFFFFFFFF8155943DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_09 = 256'h0000FFFFFFFFFFFFFFF1053C04DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0A = 256'h0000FFFFFFFFFFFFFFE09430415FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0B = 256'h0000FFFFFFFFFFFFFFE22A32B417FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0C = 256'h0000FFFFFFFFFFFFFFCA9DE25247FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0D = 256'h0000FFFFFFFFFFFFFF885DE42028B3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0E = 256'h0000FFFFFFFFFFFFFF8023C5259D6BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_0F = 256'h0000FFFFFFFFFFFFFF819AAA22003B2FFBD5D05FFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_10 = 256'h0000FFFFFFFFFFFFFEA086A850441BBCA03F3BFB6ABBBF81FFFFFFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_11 = 256'h0000FFFFFFFFFFFFFE22438054453BB8C0002120422B55AF7FF6FFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_12 = 256'h0000FFFFFFFFFFFFFE414344481466704CA525168A004102088B3FFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_13 = 256'h0000FFFFFFFFFFFFF8644B11C8003672102622D9A2C9404200465FFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_14 = 256'h0000FFFFFFFFFFFFF949D6019208EFB014DCA45D4D42A4E61313DFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_15 = 256'h0000FFFFFFFFFFFFF14D1E498912EB614D5ACADF5AB13460DA039FFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_16 = 256'h0000FFFFFFFFFFFFE41A1A435224CAE054D1322224D957D92A03AFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_17 = 256'h0000FFFFFFFFFFFFEA1A74414404BBE092DADDAFE336FB026281DFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_18 = 256'h0000FFFFFFFFFFFFCA20FA020045FCE99AFAB6B3965D2E5DB220AFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_19 = 256'h0000FFFFFFFFFFFF825CBC8265C15361D4FA2E5A2DAF72D9A248B7FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_1A = 256'h0000FFFFFFFFFFFF8049F90A112979411D345BE2D1FDA5235261BFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_1B = 256'h0000FFFFFFFFFFFF0849A1524A23D1412D5AD54D2DBD2AA5B620DFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_1C = 256'h0000FFFFFFFFFFFF31A2CA21140374831245EE053DB2D9A31A20FFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_1D = 256'h0000FFFFFFFFFFFEF0DFC21080237F44482D66DBA4DBB5B45C216BFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_1E = 256'h0000FFFFFFFFFFFCC1AB82414583E3C28DBA5DA52BB3D7AEAEA84BFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_1F = 256'h0000FFFFFFFFFFF8414DA3035025FD819DACD5DDDA35CDCB124225FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_20 = 256'h0000FFFFFFFFFFE9A54B2591B40FE7802C6ADD63DBDC1DBE62582DFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_21 = 256'h0000FFFFFFFFFFF481174DA4402EDE822DB474574D662265DA525AFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_22 = 256'h0000FFFFFFFFFFE21317024C024CD5921BB4D225E63275DCAD095AFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_23 = 256'h0000FFFFFFFFFFC91A323504901CED0125823AC55B5C5DDAED5124FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_24 = 256'h0000FFFFFFFFFFCA12142082A81DAB02D219F7CB0182E35A2D281EFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_25 = 256'h0000FFFFFFFFFF9A5A3D424A221DCF025BAC725AB526ABA7AD200D7FFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_26 = 256'h0000FFFFFFFFFE0C9AD8A5D58037AE24DD49D5EAEAA1D3DA5F10877FFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_27 = 256'h0000FFFFFFFFFC32A530A426253BAE722552D9B1AA22ACBC2A2009FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_28 = 256'h0000FFFFFFFFFF3145F020A10273556B7A004B4883C53033685E8DFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_29 = 256'h0000FFFFFFFFFE80E5B4A12010BF1BFFDF56FD75DAA9B0011200223FFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_2A = 256'h0000FFFFFFFFFFF9FEB848D49577B604082040FBBFF9FBB7DFE65FBFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_2B = 256'h0000FFFFFFFFFFF8FFDB22E620FEFC8CD445123FA821ED003C2DF3DFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_2C = 256'h0000FFFFFFFFFFBCFFEDA51C54FE5C5DA642B02BD922E448188406DFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_2D = 256'h0000FFFFFFFFFFFF7FFAD55C58E78D1AB405367FB92B6C415010837FFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_2E = 256'h0000FFFFFFFFFFFF3FFF7454196C2C558C1544277C35DC0234D183EFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_2F = 256'h0000FFFFFFFFFFFF9FFFBF08A1DC29CC041D243BEC3BF421580AC1BFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_30 = 256'h0000FFFFFFFFFFFFAFFFF2C443DAEB913E1D243B3F75A44220201ADFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_31 = 256'h0000FFFFFFFFFFFBEFFFFFF013DEF9ECA61AB43F6FFB4280402029B7FFFFFFFF;
defparam dpb_inst_0.INIT_RAM_32 = 256'h0000FFFFFFFFFFFFF7FFFFAC03FD9D5F4A15F7A37FF67ECD08AA2AF7FFFFFFFF;
defparam dpb_inst_0.INIT_RAM_33 = 256'h0000FFFFFFFFFFFEF3FFFFFFC3DB4424AE025D335C1EA210484A41DBFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_34 = 256'h0000FFFFFFFFFFFF7DFFFFFBF73A3B62CE1ABD5FA0426A0A0C4C90FFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_35 = 256'h0000FFFFFFFFFFFFFCFFFFFF7F75D16BAC2C423BE84A22450424587FFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_36 = 256'h0000FFFFFFFFFFFFFE7FFFFFEF7BF55F984A5A2FF40B7E922514A0EFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_37 = 256'h0000FFFFFFFFFFFFFF3FFFFFE777E81AA8244A3FF48DD7019408142DFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_38 = 256'h0000FFFFFFFFFFFFFF9FFFFFFEFF7FFFFFFFFDBFFA0BED8D2411B03DFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_39 = 256'h0000FFFFFFFFFFFFF7CFFFFFFFFFFFE9105FFFDEBF7FEFF7F6E64935FFFFFFFF;
defparam dpb_inst_0.INIT_RAM_3A = 256'h0000FFFFFFFFFFFFFBE7FFFFFFFFFFFFFFFFFFFFFFFFFE42FDDBBEEDFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_3B = 256'h0000FFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDBFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_3C = 256'h0000FFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF5FFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_3D = 256'h0000FFFFFFFFFFFFFFF67FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_3E = 256'h0000FFFFFFFFFFFFFFBE7FDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFF;
defparam dpb_inst_0.INIT_RAM_3F = 256'h0000FFFFFFFFFFFFFFDF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DPB dpb_inst_1 (
    .DOA({dpb_inst_1_douta_w[14:0],dpb_inst_1_douta[1]}),
    .DOB({dpb_inst_1_doutb_w[14:0],dpb_inst_1_doutb[1]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[1]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[1]})
);

defparam dpb_inst_1.READ_MODE0 = 1'b0;
defparam dpb_inst_1.READ_MODE1 = 1'b1;
defparam dpb_inst_1.WRITE_MODE0 = 2'b00;
defparam dpb_inst_1.WRITE_MODE1 = 2'b00;
defparam dpb_inst_1.BIT_WIDTH_0 = 1;
defparam dpb_inst_1.BIT_WIDTH_1 = 1;
defparam dpb_inst_1.BLK_SEL_0 = 3'b000;
defparam dpb_inst_1.BLK_SEL_1 = 3'b000;
defparam dpb_inst_1.RESET_MODE = "SYNC";
defparam dpb_inst_1.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFF92BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFE02F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFA125DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFFA202BB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_06 = 256'h0000FFFFFFFFFFFFFFFA22D677FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_07 = 256'h0000FFFFFFFFFFFFFFFC405C9CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_08 = 256'h0000FFFFFFFFFFFFFFFC043C16FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_09 = 256'h0000FFFFFFFFFFFFFFF8815AD1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0A = 256'h0000FFFFFFFFFFFFFFF21BF93A7BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0B = 256'h0000FFFFFFFFFFFFFFE015F2411EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0C = 256'h0000FFFFFFFFFFFFFFC822E201A5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0D = 256'h0000FFFFFFFFFFFFFFC440E3D1A3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0E = 256'h0000FFFFFFFFFFFFFF9CD9E082447AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_0F = 256'h0000FFFFFFFFFFFFFF58EBCD2D2C2BF77FBE2BFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_10 = 256'h0000FFFFFFFFFFFFFE19A3CA4160BD6C05EDED3FBFEEE45FFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_11 = 256'h0000FFFFFFFFFFFFFD51ADA84A81AE708829000815BDFEFBF55DFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_12 = 256'h0000FFFFFFFFFFFFFC229D11C092375A1A54428021120840445EBFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_13 = 256'h0000FFFFFFFFFFFFF9039E488691D5B81A5058044A242D004863DFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_14 = 256'h0000FFFFFFFFFFFFF90A1E7119866C7122433102BABA9210EA005FFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_15 = 256'h0000FFFFFFFFFFFFF302D42200CC2CF024453CFBA25BD31A0512DFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_16 = 256'h0000FFFFFFFFFFFFD3056D6150A06D604A5CDBDDBB66F862C190DFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_17 = 256'h0000FFFFFFFFFFFFC50259422222D868995B22445EDB25F5DC142FFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_18 = 256'h0000FFFFFFFFFFFFC51A59D641209A60A546DDAAF9E3E350498167FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_19 = 256'h0000FFFFFFFFFFFF9821D0545401BDA01A4DB32DE6659E5C3941AFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_1A = 256'h0000FFFFFFFFFFFF1C2AA285201DBFE1A5D5AA1A7E225DDDAA00C7FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_1B = 256'h0000FFFFFFFFFFFF2925D1012D81BBE2C2AD3AAAD272E55A914827FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_1C = 256'h0000FFFFFFFFFFFE585B6212921BBBE0DDB631F5C25E36DCE5D043FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_1D = 256'h0000FFFFFFFFFFFC2A42D540045361C327D5394C5A6DBA6B52586BFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_1E = 256'h0000FFFFFFFFFFFC2845E921A206B68064CB62D2D42C5AA5581075FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_1F = 256'h0000FFFFFFFFFFF9A2268D61B8DE66C042532A2225DA243DE920BBFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_20 = 256'h0000FFFFFFFFFFF0025F1CC06086F5A623AB2599AC23C2C319895AFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_21 = 256'h0000FFFFFFFFFFF24ADE14903D0DE394C2D35B54B7B9BF9E5D883DFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_22 = 256'h0000FFFFFFFFFFE48CBE9D0041CEEF0444566DF659DD5663ECE00EFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_23 = 256'h0000FFFFFFFFFFC505DD1A5A4C0FD7009A7DCE7ACAE325AE25081AFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_24 = 256'h0000FFFFFFFFFF8C15FD3A414A1BDD200DAE483DFC7A6DAFC25005FFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_25 = 256'h0000FFFFFFFFFF8445D83C0C183FAA01044B8BA5DBBB5A5A5D514D7FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_26 = 256'h0000FFFFFFFFFC2062EA50E54339DE024222222B4D3E5D2DACA01D7FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_27 = 256'h0000FFFFFFFFFC1015B45D7055BFDD3DAA18069C4FFCA287A5C80E7FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_28 = 256'h0000FFFFFFFFFE5019B5DA48813F3ED7420220A668224BD9861C0DBFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_29 = 256'h0000FFFFFFFFFE455BF06A5AA1736DDEEDFB6FBF6DEE0810000167BFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_2A = 256'h0000FFFFFFFFFEFBFDD2B4A04A7E3151450D06ADEDDE2EDAA939A5DFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_2B = 256'h0000FFFFFFFFFF79FF6E2CB9547654625610C83DF83EA005C2CB5F3FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_2C = 256'h0000FFFFFFFFFFFE7FEF899610763542221A4E7FE93FDC251422435FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_2D = 256'h0000FFFFFFFFFFBE7FFFF14409FC60D44612D15DEC35B22C18AA55DFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_2E = 256'h0000FFFFFFFFFFEF3FFFFA5141DFB922E61AB535E9B7A244102441AFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_2F = 256'h0000FFFFFFFFFFFF5FFFDF1411EFFD67D603826D2416DA14016813EFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_30 = 256'h0000FFFFFFFFFFF7CFFFFFE691BB54CEC413B23FC7B55E811C89C16FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_31 = 256'h0000FFFFFFFFFFFFE7FFFFB581B99A226A2C4537AF75A44A1C3A81D7FFFFFFFF;
defparam dpb_inst_1.INIT_RAM_32 = 256'h0000FFFFFFFFFFFFE3FFFFFEA3D2E2500D39201DA771A200A81141DBFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_33 = 256'h0000FFFFFFFFFFFFFBFFFFE7073DBBDAD53DA43DA805BA820C2240EFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_34 = 256'h0000FFFFFFFFFFFFF9FFFFF9A7BBE5BD241A443DFD592AA0A424495BFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_35 = 256'h0000FFFFFFFFFFFFBEFFFFFFDFBBFD5DD413A43EAC99ED10DA1D04DBFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_36 = 256'h0000FFFFFFFFFFFFDF7FFFFFBF6DF4A1EE2BA23769DDD24A9C525455FFFFFFFF;
defparam dpb_inst_1.INIT_RAM_37 = 256'h0000FFFFFFFFFFFFDF3FFFFFFF6D73EDA619243FF48BFAD42E5348FDFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_38 = 256'h0000FFFFFFFFFFFFFF9FFFFFFE67BF7FFFBF7FFFF9FDFE20962C4E36FFFFFFFF;
defparam dpb_inst_1.INIT_RAM_39 = 256'h0000FFFFFFFFFFFFFFCFFFFFFFFFFA02FFFFFFFFF7DB7D7F5BB0007FFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_3A = 256'h0000FFFFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFA35FFFFFEFBFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_3B = 256'h0000FFFFFFFFFFFFFDF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEEFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_3C = 256'h0000FFFFFFFFFFFFFEFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD7FFFFFFFF;
defparam dpb_inst_1.INIT_RAM_3D = 256'h0000FFFFFFFFFFFFFF7AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEDFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_3E = 256'h0000FFFFFFFFFFFFFFBF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_1.INIT_RAM_3F = 256'h0000FFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFF;

DPB dpb_inst_2 (
    .DOA({dpb_inst_2_douta_w[14:0],dpb_inst_2_douta[2]}),
    .DOB({dpb_inst_2_doutb_w[14:0],dpb_inst_2_doutb[2]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[2]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[2]})
);

defparam dpb_inst_2.READ_MODE0 = 1'b0;
defparam dpb_inst_2.READ_MODE1 = 1'b1;
defparam dpb_inst_2.WRITE_MODE0 = 2'b00;
defparam dpb_inst_2.WRITE_MODE1 = 2'b00;
defparam dpb_inst_2.BIT_WIDTH_0 = 1;
defparam dpb_inst_2.BIT_WIDTH_1 = 1;
defparam dpb_inst_2.BLK_SEL_0 = 3'b000;
defparam dpb_inst_2.BLK_SEL_1 = 3'b000;
defparam dpb_inst_2.RESET_MODE = "SYNC";
defparam dpb_inst_2.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFF097FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFF2A5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFD1AB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFFC22CDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_06 = 256'h0000FFFFFFFFFFFFFFF4444A5BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_07 = 256'h0000FFFFFFFFFFFFFFF8271E4FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_08 = 256'h0000FFFFFFFFFFFFFFF8A39A87BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_09 = 256'h0000FFFFFFFFFFFFFFF81D3829BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0A = 256'h0000FFFFFFFFFFFFFFF10839806FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0B = 256'h0000FFFFFFFFFFFFFFE6042950AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0C = 256'h0000FFFFFFFFFFFFFFC554B5D4877FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0D = 256'h0000FFFFFFFFFFFFFFC83AD00031FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0E = 256'h0000FFFFFFFFFFFFFF804B6A15147CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_0F = 256'h0000FFFFFFFFFFFFFF0002C460215D3DB6D1FFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_10 = 256'h0000FFFFFFFFFFFFFE2055846242BB347BB7BFEFED3211FFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_11 = 256'h0000FFFFFFFFFFFFFE404522C43A33394500248514EFEBBDBFEBFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_12 = 256'h0000FFFFFFFFFFFFFE23AF90542033B02A01202A8008240400ADBFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_13 = 256'h0000FFFFFFFFFFFFFCA84F20818876E0050B02AA2999A0C804225FFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_14 = 256'h0000FFFFFFFFFFFFF8C5EB00AA0267B8323C8DA9E844A9260B975FFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_15 = 256'h0000FFFFFFFFFFFFF18D3E418864EF50512246545D6604C5B2055FFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_16 = 256'h0000FFFFFFFFFFFFE2933C0B1A40DDB894022C2A4ABB579DBC022FFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_17 = 256'h0000FFFFFFFFFFFFE2AD7C4B011CDFE04D4EBDF3256DDC34C283EFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_18 = 256'h0000FFFFFFFFFFFFD4466C0320D8DD6012322A5B4E3D5D9FA4499FFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_19 = 256'h0000FFFFFFFFFFFFCC24F9024241D9E145B6BDDE11DA65A3E580D7FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_1A = 256'h0000FFFFFFFFFFFFA841F1140821D1C2541A65DF52BDA272B5A177FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_1B = 256'h0000FFFFFFFFFFFF20917580D112BAC83D22E5D52DDD3BDA7922D7FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_1C = 256'h0000FFFFFFFFFFFE2109E14002CAB64A22D5DE9A3DA1D95B14227BFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_1D = 256'h0000FFFFFFFFFFFE400B42119153BF409A2EA5A74F26CBBD5D2157FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_1E = 256'h0000FFFFFFFFFFFAC1568694260373C3122D5D5B6BB32BB5AEA45BFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_1F = 256'h0000FFFFFFFFFFFC419FC28AA2677B812DAAF5DDDA27B3CA55D825FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_20 = 256'h0000FFFFFFFFFFF98103A240A0465F819956BA6EE3D4BEBDEAA82BFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_21 = 256'h0000FFFFFFFFFFE1021349500466DE82225DDD5FDC5692E5ACE00AFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_22 = 256'h0000FFFFFFFFFFF2029621A4200E538339D95215A633995E2A1832FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_23 = 256'h0000FFFFFFFFFFC4223CA50D001CCF826542A59B2D3DDA65D5E44EFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_24 = 256'h0000FFFFFFFFFF855A2C4A01259DAF0162A1B7C59B36B2A57B0A3A7FFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_25 = 256'h0000FFFFFFFFFFCA225C4530861DDF01B2ACF57A5E64ADADA6800D7FFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_26 = 256'h0000FFFFFFFFFD1C1CB85A41081FAB002999DDAD22A5A3DAD618057FFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_27 = 256'h0000FFFFFFFFFA14EAF9402A21359E0F05CAD262209F5A705421057FFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_28 = 256'h0000FFFFFFFFFF19CCF04A01403BDD2800255A5126D9342CB98C06FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_29 = 256'h0000FFFFFFFFFE32A1B90900313F33ED775FF7D5B650AA8AA00085BFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2A = 256'h0000FFFFFFFFFEF9FEF881DD0A77DE0A20A2DBFF7EFBBB7DE7CE6ABFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2B = 256'h0000FFFFFFFFFFFCFFBD10CC00DFBD0A240A057FD823FAD81F75DDDFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2C = 256'h0000FFFFFFFFFFF9FFEBC6A4A8FDF915B605223EB8226100A4A007DFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2D = 256'h0000FFFFFFFFFFFE7FFB611AA4EE2D23351D5C3FF815ED012245036FFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2E = 256'h0000FFFFFFFFFFFF3FFEBC4C98ECEDBE1287523FD814FA21109222FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_2F = 256'h0000FFFFFFFFFFEF9FFFDB9191DD98996D3C1E36DC336C41580541BFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_30 = 256'h0000FFFFFFFFFFF7DFFFF68049DCFB715E1CD53FFFF4A4C8404623B7FFFFFFFF;
defparam dpb_inst_2.INIT_RAM_31 = 256'h0000FFFFFFFFFFFFCFFFFCF023DEEBDAAD03A23FE7F2BAA4408628FFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_32 = 256'h0000FFFFFFFFFFFBF7FFFF5C23BDBDD16C0ED523EF7DEC944A69106FFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_33 = 256'h0000FFFFFFFFFFFEF3FFFFEFA3D5E46E4C12AB5BCC1AE640D02914F7FFFFFFFF;
defparam dpb_inst_2.INIT_RAM_34 = 256'h0000FFFFFFFFFFFFFBFFFFFBE7DA5AA6BD25A91F4C0AEA4A1C2120EFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_35 = 256'h0000FFFFFFFFFFFFFCFFFFFEFFB2C2CA5A2CD33FF41A12842C80E0ADFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_36 = 256'h0000FFFFFFFFFFFFFE7FFFFFDFB563BEAC14593BBC0AD944420920FDFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_37 = 256'h0000FFFFFFFFFFFFFF3FFFFFEF67EC92DC469236BA0D7E02840C286DFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_38 = 256'h0000FFFFFFFFFFFFEFBFFFFFFEFFFFFFFFFB80BFF7BBB7044C02403DFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_39 = 256'h0000FFFFFFFFFFFFF7CFFFFFFFFD21DFFFFFFFFFFFFFFFF5FA912A5AFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3A = 256'h0000FFFFFFFFFFFFFBEFFFFF7FFFFFFFBFFFFFFFFFF017F6BDBDFBEBFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3B = 256'h0000FFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3C = 256'h0000FFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3D = 256'h0000FFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3E = 256'h0000FFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEBFFFFFFFFF;
defparam dpb_inst_2.INIT_RAM_3F = 256'h0000FFFFFFFFFFFFFFDFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFFF;

DPB dpb_inst_3 (
    .DOA({dpb_inst_3_douta_w[14:0],dpb_inst_3_douta[3]}),
    .DOB({dpb_inst_3_doutb_w[14:0],dpb_inst_3_doutb[3]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[3]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[3]})
);

defparam dpb_inst_3.READ_MODE0 = 1'b0;
defparam dpb_inst_3.READ_MODE1 = 1'b1;
defparam dpb_inst_3.WRITE_MODE0 = 2'b00;
defparam dpb_inst_3.WRITE_MODE1 = 2'b00;
defparam dpb_inst_3.BIT_WIDTH_0 = 1;
defparam dpb_inst_3.BIT_WIDTH_1 = 1;
defparam dpb_inst_3.BLK_SEL_0 = 3'b000;
defparam dpb_inst_3.BLK_SEL_1 = 3'b000;
defparam dpb_inst_3.RESET_MODE = "SYNC";
defparam dpb_inst_3.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFFBA7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFE847FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFD28DDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFFE1057AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_06 = 256'h0000FFFFFFFFFFFFFFFE211E7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_07 = 256'h0000FFFFFFFFFFFFFFF041941AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_08 = 256'h0000FFFFFFFFFFFFFFFC8C5C22FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_09 = 256'h0000FFFFFFFFFFFFFFF982AA04EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0A = 256'h0000FFFFFFFFFFFFFFF187D0427FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0B = 256'h0000FFFFFFFFFFFFFFE139F00A37FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0C = 256'h0000FFFFFFFFFFFFFFE02AE0215FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0D = 256'h0000FFFFFFFFFFFFFF8245ECB1A16FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0E = 256'h0000FFFFFFFFFFFFFFCC51C542046DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_0F = 256'h0000FFFFFFFFFFFFFF2CDBC228103B77DD3FFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_10 = 256'h0000FFFFFFFFFFFFFF09A2D920412BFFFFFBEBF777FDDFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_11 = 256'h0000FFFFFFFFFFFFFE19A39856895BF100150040FFBDFFEEFA2BFFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_12 = 256'h0000FFFFFFFFFFFFFC50469841117ED839000400494100202EF7FFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_13 = 256'h0000FFFFFFFFFFFFFA474B19C4C6563014A4DCA3A442420240375FFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_14 = 256'h0000FFFFFFFFFFFFFD021E39901276E4120370AA4BA2545106035FFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_15 = 256'h0000FFFFFFFFFFFFF0849D2984022CF04AD53305025A7A584923BFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_16 = 256'h0000FFFFFFFFFFFFF20C3D612D00CCE423B5A5E5A6AD98E04123DFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_17 = 256'h0000FFFFFFFFFFFFCC143D231402D8612231DA1D9132E35269012FFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_18 = 256'h0000FFFFFFFFFFFFC521B8C25041BBD1A9DDADADF364A4605301EFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_19 = 256'h0000FFFFFFFFFFFF821AD9942D053D61124AC667EF2DB27D78495FFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_1A = 256'h0000FFFFFFFFFFFF041DB88640993D6103E5BAA1EDD5BB5AE04897FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_1B = 256'h0000FFFFFFFFFFFF1C4BD0940883B54282DD5A2FD562A42B9580B7FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_1C = 256'h0000FFFFFFFFFFFE54A755100029F5C15C35626DC2BEE6ADE1109FFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_1D = 256'h0000FFFFFFFFFFFE3163E1888806E1C2A5D3DAD9B5F12E4DA8C85BFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_1E = 256'h0000FFFFFFFFFFFC528BD240C2177A949BE162AA54DDA4DA51502BFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_1F = 256'h0000FFFFFFFFFFF8A2C52C42D823E6C2925B1A5246B9DD6B58003BFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_20 = 256'h0000FFFFFFFFFFFAA2DD0D12720FE284AF9DE5A23CBA42D6AC902DFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_21 = 256'h0000FFFFFFFFFFF08D5F86AC649EEB855BA2ABE6E331EA3AA2123BFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_22 = 256'h0000FFFFFFFFFFE2055E1C1A61CBEF0086275DFAD1DC6DF5EDA11DFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_23 = 256'h0000FFFFFFFFFFE31AAE1208AA0EF311193AF2CAE792A55AAA1022FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_24 = 256'h0000FFFFFFFFFFC8056D2A11101DEB082D5ECC7C4EDBAAB504A00DFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_25 = 256'h0000FFFFFFFFFF145D6920184135AD2085569A9FE3BB56A6DC78177FFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_26 = 256'h0000FFFFFFFFFE2042E948A3B5BDAE0184AA0562BDB45DAE2DC12F7FFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_27 = 256'h0000FFFFFFFFFF1005509A50623B6A03D2291D359A65C59FDAD89FBFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_28 = 256'h0000FFFFFFFFFC602B3CA5C5183F1F8000110B4A902642A246688ABFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_29 = 256'h0000FFFFFFFFFFC1BAE1E498DDF74AF7DDB55DFF920404A414C5C6FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2A = 256'h0000FFFFFFFFFE75FBB178C2063E324002297DDDAB6BED8E1C330B7FFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2B = 256'h0000FFFFFFFFFF79FF6E2AE5627664A25720A02B687DA825B5DD67FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2C = 256'h0000FFFFFFFFFF7CFFEF025A146E3C64CA1AD13FE93BDC5A1202855FFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2D = 256'h0000FFFFFFFFFFBE7FFBE94C28FF545DD604A23DE93B54A23010C6DFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2E = 256'h0000FFFFFFFFFFFFBFFED95041FF2040EE199D2F6C339D12B8598B6FFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_2F = 256'h0000FFFFFFFFFFFF3FFFDE1449ECEA655400A12B281FE614225292EFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_30 = 256'h0000FFFFFFFFFFFFCFFFF7A523DF215AC51A027AAE3FD402103491FFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_31 = 256'h0000FFFFFFFFFFFBEFFFFFF111D935654C3C957DBF7D4C01586089B7FFFFFFFF;
defparam dpb_inst_3.INIT_RAM_32 = 256'h0000FFFFFFFFFFFFE7FFFF7A61DAD20DAEA5251FD7725622280A89B7FFFFFFFF;
defparam dpb_inst_3.INIT_RAM_33 = 256'h0000FFFFFFFFFFFFFBFFFFDB03BA3B23AC1AE4242917502A1C5240BBFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_34 = 256'h0000FFFFFFFFFFFEF9FFFFFBC73D25B5CC1AAA37A19ABA014814883BFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_35 = 256'h0000FFFFFFFFFFFFFDFFFFFEBF7F7A6DAC16585D599DEA520C2A1CFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_36 = 256'h0000FFFFFFFFFFFFBEFFFFFF9F77F452DC3BA23FE4AB66028C221457FFFFFFFF;
defparam dpb_inst_3.INIT_RAM_37 = 256'h0000FFFFFFFFFFFFDF7FFFFFEF7BE27E8419EA3FF48BED522E11886DFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_38 = 256'h0000FFFFFFFFFFFFEF9FFFFFFC67DFFFFFE4543B728DFD52261114F7FFFFFFFF;
defparam dpb_inst_3.INIT_RAM_39 = 256'h0000FFFFFFFFFFFFFFAFFFFFFFE41FFFFFBFFFFFFFFDEFFF882C843FFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_3A = 256'h0000FFFFFFFFFFFFFFE7FFFFFFFFFEFFFFFFFFFF340DFEBFFFFF7EBEFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_3B = 256'h0000FFFFFFFFFFFFFDF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF41DFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_3C = 256'h0000FFFFFFFFFFFFFFF9EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_3D = 256'h0000FFFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_3E = 256'h0000FFFFFFFFFFFFFFBE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFF;
defparam dpb_inst_3.INIT_RAM_3F = 256'h0000FFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFFFFFFF;

DPB dpb_inst_4 (
    .DOA({dpb_inst_4_douta_w[11:0],dpb_inst_4_douta[3:0]}),
    .DOB({dpb_inst_4_doutb_w[11:0],dpb_inst_4_doutb[3:0]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[14],ada[13],ada[12]}),
    .BLKSELB({adb[14],adb[13],adb[12]}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[3:0]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[3:0]})
);

defparam dpb_inst_4.READ_MODE0 = 1'b0;
defparam dpb_inst_4.READ_MODE1 = 1'b1;
defparam dpb_inst_4.WRITE_MODE0 = 2'b00;
defparam dpb_inst_4.WRITE_MODE1 = 2'b00;
defparam dpb_inst_4.BIT_WIDTH_0 = 4;
defparam dpb_inst_4.BIT_WIDTH_1 = 4;
defparam dpb_inst_4.BLK_SEL_0 = 3'b100;
defparam dpb_inst_4.BLK_SEL_1 = 3'b100;
defparam dpb_inst_4.RESET_MODE = "SYNC";
defparam dpb_inst_4.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFFEFFF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_02 = 256'hFFFFFFFFFFF5FFFFF50FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_03 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFFFEDBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_06 = 256'hFFFFFFFFFFFFAFFFFF14EFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_07 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFBFFDBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_0A = 256'hFFFFFFFFFFFFF7AFFFF24DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_0B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_0C = 256'hFFFFFFFFFFFFDFFFDBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFBFFFFF50EFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_0F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_10 = 256'hFFFFFFFFFFFFFFDB7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFF6FFFFF82DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_13 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_14 = 256'hFFFFFFFFFFFFDB7DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFF7FFFF6B0EFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_17 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_18 = 256'hFFFFFFD9EC8812BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFFF6FFFF24DFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1C = 256'hFFFFFA51112A1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFFAFFFF12DFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_1F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_20 = 256'hFFFDBCA88030FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFFFAFFFF58BFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFEFFFFF;
defparam dpb_inst_4.INIT_RAM_23 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_24 = 256'hFFF5657DA52FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7F;
defparam dpb_inst_4.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFFBFFFF50FFFFFFBFFFFFFFFFFFFFFFFFFFFFFF7FFFFF;
defparam dpb_inst_4.INIT_RAM_27 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_28 = 256'hFFFFFFBF57FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_29 = 256'hFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFFF2FFFF74DFFFFFFFFFFDFFFFFFFFFFFFFF7FFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2C = 256'hFFD7F7CBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2D = 256'hFFFFFFFFFFFF7FFFFFFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFFF7EFFF40DFFFFFBFFFFFBFFFFFFFFFEDFF7FFFFFFB;
defparam dpb_inst_4.INIT_RAM_2F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_30 = 256'hFEBF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_31 = 256'hDBBBB3FBBBBBBB9BBFBBB36BB3FB37737777777F7FF7E3FFFFFFFFF7FFFFBFFF;
defparam dpb_inst_4.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFF7D7DDCC9DF9BDBDADDBDDB9FCBBD9FDBB9B5;
defparam dpb_inst_4.INIT_RAM_33 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_35 = 256'hFFFBFFFB7FFFFFFFFFFFFFFFFF7F7FFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFF33FFDFB7FFFFFFFFBFFFBFFFBFFFFF;
defparam dpb_inst_4.INIT_RAM_37 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_4.INIT_RAM_3F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DPB dpb_inst_5 (
    .DOA({dpb_inst_5_douta_w[14:0],dpb_inst_5_douta[4]}),
    .DOB({dpb_inst_5_doutb_w[14:0],dpb_inst_5_doutb[4]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[4]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[4]})
);

defparam dpb_inst_5.READ_MODE0 = 1'b0;
defparam dpb_inst_5.READ_MODE1 = 1'b1;
defparam dpb_inst_5.WRITE_MODE0 = 2'b00;
defparam dpb_inst_5.WRITE_MODE1 = 2'b00;
defparam dpb_inst_5.BIT_WIDTH_0 = 1;
defparam dpb_inst_5.BIT_WIDTH_1 = 1;
defparam dpb_inst_5.BLK_SEL_0 = 3'b000;
defparam dpb_inst_5.BLK_SEL_1 = 3'b000;
defparam dpb_inst_5.RESET_MODE = "SYNC";
defparam dpb_inst_5.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFFDDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFE021FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFE067FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFFF420DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_06 = 256'h0000FFFFFFFFFFFFFFF8824D6BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_07 = 256'h0000FFFFFFFFFFFFFFFA049F0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_08 = 256'h0000FFFFFFFFFFFFFFF841AD8F7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_09 = 256'h0000FFFFFFFFFFFFFFF88D7DD3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0A = 256'h0000FFFFFFFFFFFFFFF02879386FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0B = 256'h0000FFFFFFFFFFFFFFE00AB5A03EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0C = 256'h0000FFFFFFFFFFFFFFC222719185FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0D = 256'h0000FFFFFFFFFFFFFFC458E24533FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0E = 256'h0000FFFFFFFFFFFFFF002EE22212F5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_0F = 256'h0000FFFFFFFFFFFFFF90A16922642F5BE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_10 = 256'h0000FFFFFFFFFFFFFF201B44522DBA5EDFFEBF5DDA7FFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_11 = 256'h0000FFFFFFFFFFFFFE42D78448443E3B4480941DAAEEDAFB27C7FFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_12 = 256'h0000FFFFFFFFFFFFFE031782C04016B26014010800088201935A3FFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_13 = 256'h0000FFFFFFFFFFFFFC22A720A9037BF9112202145324100002153FFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_14 = 256'h0000FFFFFFFFFFFFF0D54B848A825C7019BD0A4DA45A432C93C5DFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_15 = 256'h0000FFFFFFFFFFFFFAA226210160EE58244BDCB2D95B05252402CFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_16 = 256'h0000FFFFFFFFFFFFF143948311896FA05852D216596A252DA601AFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_17 = 256'h0000FFFFFFFFFFFFE3015CC1825C5DE0ADCC2DA5FFDD395AC4A1AFFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_18 = 256'h0000FFFFFFFFFFFFE4145A222920CC608A56E2E43D3B5B9518802FFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_19 = 256'h0000FFFFFFFFFFFFDC4270868415D9A2D9A535953ED5DB840601A7FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_1A = 256'h0000FFFFFFFFFFFF9840D52404A3B3C1BC1A5ABED26ADDEE3A01B7FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_1B = 256'h0000FFFFFFFFFFFE80A4E200CD0373C15D2225D02BBDDBBC5AA0D7FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_1C = 256'h0000FFFFFFFFFFFE3091E2A8902B33428BDE5B523CA15AA61EA0E3FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_1D = 256'h0000FFFFFFFFFFFC512EAA2685A37E425AAC6D4EFD1AA3B2D6206BFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_1E = 256'h0000FFFFFFFFFFFC0066C52011136FC1543F5AA54A22BB5A9A10CBFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_1F = 256'h0000FFFFFFFFFFFC0027830A20EE7390ADA4E5CD3555E2ADAEE92DFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_20 = 256'h0000FFFFFFFFFFF0002FA28988067FC204E45A5DDEABBA2B424955FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_21 = 256'h0000FFFFFFFFFFF2411D5A41C8E66FC40ABEF6755DDA1DCDFDD82DFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_22 = 256'h0000FFFFFFFFFFF1909343C1280DD3A2D5B962451E63975E54182EFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_23 = 256'h0000FFFFFFFFFFC402565DAA00AA9D0247CE9AE52D7A5B2E5C481AFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_24 = 256'h0000FFFFFFFFFF8A2A5429854A1D9F0125EA7383E126DDDDFA49167FFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_25 = 256'h0000FFFFFFFFFF8A023C5E488C1BD70275246FEA2C955DDA260019FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_26 = 256'h0000FFFFFFFFFE1E3A3C2644101BD7107145F29FCAB3A2F5D228057FFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_27 = 256'h0000FFFFFFFFFF3862BC4938213F9F4714A4D592A59272A42E40027FFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_28 = 256'h0000FFFFFFFFFE19C5E25805013BB5010194A4156D513A4D51080D7FFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_29 = 256'h0000FFFFFFFFFE324B781120467B373D65DBF6A02022D2516000133FFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_2A = 256'h0000FFFFFFFFFEF3FFD80AD41277DC015D6FAF7FFFFEAEF5E38007BFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_2B = 256'h0000FFFFFFFFFFF9FF7558E90277B215040A047FBFA6DFDADA22BA5FFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_2C = 256'h0000FFFFFFFFFFFAFFB79A25A0F6ED1226055C3DF927790488504FAFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_2D = 256'h0000FFFFFFFFFFDE7FF7C2A284ED292224965E3F6915EC1918AA05BFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_2E = 256'h0000FFFFFFFFFFDE7FFFF48D18ECDD5F1484A537F83EE448000223AFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_2F = 256'h0000FFFFFFFFFFEF9FFFBF5211DDAD9E86227A3DEDB55441100843DFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_30 = 256'h0000FFFFFFFFFFF79FFFFFC861E8DCC92E05E52FE7F2F48198A242D7FFFFFFFF;
defparam dpb_inst_5.INIT_RAM_31 = 256'h0000FFFFFFFFFFFFEFFFFDE983DDDA55AE02A32FEE33A4C8083281DFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_32 = 256'h0000FFFFFFFFFFFFF7FFFFBC83BDD592C415A42FEF7BE0420C2441EFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_33 = 256'h0000FFFFFFFFFFFFF3FFFFCFA3BBD5DCD65C153BACFDFE00180D18DBFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_34 = 256'h0000FFFFFFFFFFFF79FFFFFBC3BBB4DA6E1C553FDC89E644082289EFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_35 = 256'h0000FFFFFFFFFFFF7CFFFFFFDFB2A296DC19AB3FAC8212022C2440ABFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_36 = 256'h0000FFFFFFFFFFFFFC7FFFFFFFB6B7AD4A0C5A3BF48999506A19D0FDFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_37 = 256'h0000FFFFFFFFFFFFFF3FFFFFDF6EF352DC1A443BFC09BE24A4842A77FFFFFFFF;
defparam dpb_inst_5.INIT_RAM_38 = 256'h0000FFFFFFFFFFFFFF3FFFFFFA7DFF7FFD11003FFE1BFF008A1AAA5DFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_39 = 256'h0000FFFFFFFFFFFFF7CFFFFFFF89FFFFFFFFFFDEFEBFFB600284525EFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_3A = 256'h0000FFFFFFFFFFFFFFCFFFFFFFFFFFFFFFFFED2085FBEBDDFFDFDFEFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_3B = 256'h0000FFFFFFFFFFFFFFF7DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF1DE7FFFFFFFF;
defparam dpb_inst_5.INIT_RAM_3C = 256'h0000FFFFFFFFFFFFFEFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDF7FFFFFFFF;
defparam dpb_inst_5.INIT_RAM_3D = 256'h0000FFFFFFFFFFFFFFFAFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF6FFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_3E = 256'h0000FFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFF;
defparam dpb_inst_5.INIT_RAM_3F = 256'h0000FFFFFFFFFFFFFFDF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DPB dpb_inst_6 (
    .DOA({dpb_inst_6_douta_w[14:0],dpb_inst_6_douta[5]}),
    .DOB({dpb_inst_6_doutb_w[14:0],dpb_inst_6_doutb[5]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[5]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[5]})
);

defparam dpb_inst_6.READ_MODE0 = 1'b0;
defparam dpb_inst_6.READ_MODE1 = 1'b1;
defparam dpb_inst_6.WRITE_MODE0 = 2'b00;
defparam dpb_inst_6.WRITE_MODE1 = 2'b00;
defparam dpb_inst_6.BIT_WIDTH_0 = 1;
defparam dpb_inst_6.BIT_WIDTH_1 = 1;
defparam dpb_inst_6.BLK_SEL_0 = 3'b000;
defparam dpb_inst_6.BLK_SEL_1 = 3'b000;
defparam dpb_inst_6.RESET_MODE = "SYNC";
defparam dpb_inst_6.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFF296FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFD1157FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFFE19E6BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_06 = 256'h0000FFFFFFFFFFFFFFF8112EBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_07 = 256'h0000FFFFFFFFFFFFFFF0A154B2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_08 = 256'h0000FFFFFFFFFFFFFFFD0A34437FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_09 = 256'h0000FFFFFFFFFFFFFFF84018016FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0A = 256'h0000FFFFFFFFFFFFFFF9863985B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0B = 256'h0000FFFFFFFFFFFFFFE524F04917FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0C = 256'h0000FFFFFFFFFFFFFFE81DDA24CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0D = 256'h0000FFFFFFFFFFFFFFD0226931D3BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0E = 256'h0000FFFFFFFFFFFFFFCA51C98508BBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_0F = 256'h0000FFFFFFFFFFFFFF089BC4A121333C3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_10 = 256'h0000FFFFFFFFFFFFFF99A3C26A143FBB76BFFBF7E5FFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_11 = 256'h0000FFFFFFFFFFFFFE2021D8C40033F1004445EEFBFF6F57B83FFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_12 = 256'h0000FFFFFFFFFFFFFE34E558404976F0348240401024285EFFFFFFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_13 = 256'h0000FFFFFFFFFFFFFD025B92AC8026B01490A16914D10922004FDFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_14 = 256'h0000FFFFFFFFFFFFF8059E22C03067510C45D2341185388220825FFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_15 = 256'h0000FFFFFFFFFFFFF20DBD519D906774112407450571A5849A223FFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_16 = 256'h0000FFFFFFFFFFFFF30C7E515404E4E04D9439D9ADA5BC61D120DFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_17 = 256'h0000FFFFFFFFFFFFE49B344A4040DAA04023A2DA0022DD255A04CFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_18 = 256'h0000FFFFFFFFFFFFC539FC8B22C9BBD0A5533A5B9FECA475C621AFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_19 = 256'h0000FFFFFFFFFFFF8535BA904895DFE10E7AB4EFD5AC5C7371C4DFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_1A = 256'h0000FFFFFFFFFFFF9A15F0844291DAE003E5AA655D5A265161A0EFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_1B = 256'h0000FFFFFFFFFFFF3C1371469001B9C022DBFA6FD6522EC7D048B7FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_1C = 256'h0000FFFFFFFFFFFF184B31040251FDC024A52D4BC3BFADFDE150BFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_1D = 256'h0000FFFFFFFFFFFE49A3E581F20363C00AB356F742EDBE4E6998ABFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_1E = 256'h0000FFFFFFFFFFFCA2134280009762841BC4AD5ABBFAA4AFBDD873FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_1F = 256'h0000FFFFFFFFFFF9D355ADC3B0475E84925B3A35956C3D2A5820B3FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_20 = 256'h0000FFFFFFFFFFF9D3158DA2F605E582E23B65A223E4CDD4FB302DFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_21 = 256'h0000FFFFFFFFFFF905A505A0244DE50362D45B5E243DE63644415CFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_22 = 256'h0000FFFFFFFFFFE20A3F1828C40EDF041245DDB7E29CFAA32BC811FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_23 = 256'h0000FFFFFFFFFFE1953E2405204FEF2158A0ED3A9515A5B3A7A81EFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_24 = 256'h0000FFFFFFFFFFC4153E9204251DEB81A2258CFC3EB5642505202BFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_25 = 256'h0000FFFFFFFFFF8435A90530D13DDB0119DBD23BB375A42DD9980E7FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_26 = 256'h0000FFFFFFFFFE0005D0D4035A3DBA040A5A4D60665CDF565D201D7FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_27 = 256'h0000FFFFFFFFFC093DD2A4CAC23B5C00A225A85A52753AB7D9201FBFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_28 = 256'h0000FFFFFFFFFC201CB08493183F5E2020A213A2125D42B55DA40FBFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_29 = 256'h0000FFFFFFFFFE4165A45C92316F9BE2BAAD5C510ADC492D1E5B0DFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_2A = 256'h0000FFFFFFFFFE79E3E5A422847E222A45F6FFEBAEDD73AA181105BFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_2B = 256'h0000FFFFFFFFFF79FF5C45E2837E6CA0C200A177EF9B6A6B5FFFDFFFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_2C = 256'h0000FFFFFFFFFF7CFFFB0D6A107F346BA514426FD835CCA2012006FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_2D = 256'h0000FFFFFFFFFFFEFFF6D21A60EDDCCDAA09253FF83B7482A40242DFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_2E = 256'h0000FFFFFFFFFFFE3FFEF0E481EFAA21E61A50BDED23BA02B8A882FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_2F = 256'h0000FFFFFFFFFFFFBFFFEC2941EEF8A01A1BCD455817FA1452A212E7FFFFFFFF;
defparam dpb_inst_6.INIT_RAM_30 = 256'h0000FFFFFFFFFFFFAFFFE58D11BFF326A55A3275AFFD1A3A1059137FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_31 = 256'h0000FFFFFFFFFFFFCFFFF9E251DED1BA463A543FEF74D205100829F7FFFFFFFF;
defparam dpb_inst_6.INIT_RAM_32 = 256'h0000FFFFFFFFFFFBE7FFFED863DA72FADE1A5356D73D5E92A0B110B7FFFFFFFF;
defparam dpb_inst_6.INIT_RAM_33 = 256'h0000FFFFFFFFFFFDF7FFFFFE13DCDA2A6A0B421DA7F6422D882082FFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_34 = 256'h0000FFFFFFFFFFFFFBFFFFFFC7DDD3274423A23BA91A5311AD1054BBFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_35 = 256'h0000FFFFFFFFFFFFB9FFFFFEFFBDDED44546441FE499BE11802124EBFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_36 = 256'h0000FFFFFFFFFFFFBEFFFFFF3F75D0D5AC2BA55FBC4AE6090C44182FFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_37 = 256'h0000FFFFFFFFFFFFDF7FFFFFEF63E95D5545B93F629EE3014C32C05DFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_38 = 256'h0000FFFFFFFFFFFFEF1FFFFFFB67BFF54088553FE40ADD5A2C400075FFFFFFFF;
defparam dpb_inst_6.INIT_RAM_39 = 256'h0000FFFFFFFFFFFFFFDFFFFFFFD2FFFFFFFFFFFFF7DB7F905C51083BFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_3A = 256'h0000FFFFFFFFFFFFFBE7FFFFFFFFFFFFFFEBF5AFFDDEBFFF77FAF5B7FFFFFFFF;
defparam dpb_inst_6.INIT_RAM_3B = 256'h0000FFFFFFFFFFFFFDF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE0FF79FFFFFFFF;
defparam dpb_inst_6.INIT_RAM_3C = 256'h0000FFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_3D = 256'h0000FFFFFFFFFFFFFEFCDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_3E = 256'h0000FFFFFFFFFFFFFFFE7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFF;
defparam dpb_inst_6.INIT_RAM_3F = 256'h0000FFFFFFFFFFFFFFFE3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFF;

DPB dpb_inst_7 (
    .DOA({dpb_inst_7_douta_w[14:0],dpb_inst_7_douta[6]}),
    .DOB({dpb_inst_7_doutb_w[14:0],dpb_inst_7_doutb[6]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[6]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[6]})
);

defparam dpb_inst_7.READ_MODE0 = 1'b0;
defparam dpb_inst_7.READ_MODE1 = 1'b1;
defparam dpb_inst_7.WRITE_MODE0 = 2'b00;
defparam dpb_inst_7.WRITE_MODE1 = 2'b00;
defparam dpb_inst_7.BIT_WIDTH_0 = 1;
defparam dpb_inst_7.BIT_WIDTH_1 = 1;
defparam dpb_inst_7.BLK_SEL_0 = 3'b000;
defparam dpb_inst_7.BLK_SEL_1 = 3'b000;
defparam dpb_inst_7.RESET_MODE = "SYNC";
defparam dpb_inst_7.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFF863FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFE827BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFFF004BDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_06 = 256'h0000FFFFFFFFFFFFFFFC2597EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_07 = 256'h0000FFFFFFFFFFFFFFF8461E3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_08 = 256'h0000FFFFFFFFFFFFFFF8459E1FBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_09 = 256'h0000FFFFFFFFFFFFFFF90BBAD3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0A = 256'h0000FFFFFFFFFFFFFFF013B220FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0B = 256'h0000FFFFFFFFFFFFFFF21A75243DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0C = 256'h0000FFFFFFFFFFFFFFE24461D21BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0D = 256'h0000FFFFFFFFFFFFFFCA1DE54A26FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0E = 256'h0000FFFFFFFFFFFFFF804CE46080DBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_0F = 256'h0000FFFFFFFFFFFFFF802AE261403BC7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_10 = 256'h0000FFFFFFFFFFFFFE00CA9C4549336FBFEAEF544FFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_11 = 256'h0000FFFFFFFFFFFFFE119F8450213A3A11125ADBAEDBB3DAC5FFFFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_12 = 256'h0000FFFFFFFFFFFFFD431B8093852B58E0000409490105AB7DBD7FFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_13 = 256'h0000FFFFFFFFFFFFFCA14E50882B765C0A1E9502A204441010023FFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_14 = 256'h0000FFFFFFFFFFFFF9A44E90080C3DB0021229CDA4D4C22400A39FFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_15 = 256'h0000FFFFFFFFFFFFF18256448A0065A02C9BB058E4ACD4B24103DFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_16 = 256'h0000FFFFFFFFFFFFF123142322026AD0245ACE2CBE79432A9A0B4FFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_17 = 256'h0000FFFFFFFFFFFFEA44DC43022A4DF05ED8BA2ABFFD5AF4A2037FFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_18 = 256'h0000FFFFFFFFFFFFD20428A2BC00DCE8996CCDAAE3A37B92A289AFFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_19 = 256'h0000FFFFFFFFFFFFD208F8862015B0A0A14D5B77D273AB958A00E7FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_1A = 256'h0000FFFFFFFFFFFF8958B91520C9BB63AC3A6F9BA5A5D7FD9A40B7FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_1B = 256'h0000FFFFFFFFFFFF0049D9180D22BBC39D2A2B916B3DE2382B24D7FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_1C = 256'h0000FFFFFFFFFFFE2111C450401B3363BAD7A5B53CD6A2021A48C7FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_1D = 256'h0000FFFFFFFFFFFE325AC2201B03BD43A64A6F5A3D3243B524446FFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_1E = 256'h0000FFFFFFFFFFFCB1CFA2288A53FDC1CC336AEA442ADBF454045BFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_1F = 256'h0000FFFFFFFFFFFC20A782015106E3C24DAAD2A4D593DBE7AE982DFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_20 = 256'h0000FFFFFFFFFFF804CEA24A210E7E801DAD5ADDDA3A222F088275FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_21 = 256'h0000FFFFFFFFFFF0C21F9A41502EEF841E5B2DA3DBD215DDB22827FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_22 = 256'h0000FFFFFFFFFFF0499B4D92628EED82ADBC32551A73BB7DDC253EFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_23 = 256'h0000FFFFFFFFFFEA15951322105CEB810ADE52A5FAF67ACCDC4222FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_24 = 256'h0000FFFFFFFFFFCB05A42D84901ADE4059DA7A2743DA5BDDF198147FFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_25 = 256'h0000FFFFFFFFFFDA4A7C6415451EAE21C22C5DCCCC9A7BA624A815FFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_26 = 256'h0000FFFFFFFFFF1CAA7A1204221FCF216525B3BF55377555AD94077FFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_27 = 256'h0000FFFFFFFFFD2802685A70082FAE0255500BA5DA99DED42ED0067FFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_28 = 256'h0000FFFFFFFFFD5CA3D4BA0551B3AE820A59C859C9225DCA04A0857FFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_29 = 256'h0000FFFFFFFFFF3119F18040423B5EBFEFB6220CE24115D2C123063FFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_2A = 256'h0000FFFFFFFFFF33FDF051980037DD95BF5BD6BEF56B5E55210012BFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_2B = 256'h0000FFFFFFFFFFFDFFF468589277BE1A2492107EE05DBFBDE5AA6B1FFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_2C = 256'h0000FFFFFFFFFFF8FFDFA2A654E6DD04D609293EE912B410AA0C1B5FFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_2D = 256'h0000FFFFFFFFFFBC7FFBA59D1CEE2C22D515B0B6A915CA2810D183DFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_2E = 256'h0000FFFFFFFFFFFEBFFDB92C28ECA59A1C8D9E3F5835ED28144A43AFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_2F = 256'h0000FFFFFFFFFFEF5FFFBE2218EA4A40CE0A2A3B6932C509185941BFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_30 = 256'h0000FFFFFFFFFFFF9FFFFF00D9DC59F34A0DA45FEFB7DC84540441EFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_31 = 256'h0000FFFFFFFFFFF3EFFFFDE223D95BC5DC0DA276AFF25CD0DA46815FFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_32 = 256'h0000FFFFFFFFFFFFF7FFFFF891DB5D06A62DA41FEF774048184A29F7FFFFFFFF;
defparam dpb_inst_7.INIT_RAM_33 = 256'h0000FFFFFFFFFFFFF3FFFFDF03BB2DAF9C385522FFF3BE405CA6282BFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_34 = 256'h0000FFFFFFFFFFFFFBFFFFF38335AAB4BE3A3D3ECC1BF404108500EFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_35 = 256'h0000FFFFFFFFFFFFFCFFFFFFFFEA52BBBC19B537D81A424A2E1A103BFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_36 = 256'h0000FFFFFFFFFFFFFEFFFFFFEFBBF56DAA14503EE01A12422A2245F5FFFFFFFF;
defparam dpb_inst_7.INIT_RAM_37 = 256'h0000FFFFFFFFFFFFFE3FFFFFDFFE75AB9832463FFC0BFE54240A5A6BFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_38 = 256'h0000FFFFFFFFFFFFFFBFFFFFF37BF7DA2C45003EF68F7700862ADC3DFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_39 = 256'h0000FFFFFFFFFFFFEF8FFFFFFF37EFFFFFFFDBFF7DFFDE0D0014A22EFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_3A = 256'h0000FFFFFFFFFFFFFFCFFFFFFFFFFFFFFDFD0AEDFFFFFFFFBEEF5EBEFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_3B = 256'h0000FFFFFFFFFFFFFBF7FFFFFFFFFFFFFFFFFFFFFFFFFFF7521FEFFDFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_3C = 256'h0000FFFFFFFFFFFFFEFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_3D = 256'h0000FFFFFFFFFFFFFFF9FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_3E = 256'h0000FFFFFFFFFFFFFF7E7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFF;
defparam dpb_inst_7.INIT_RAM_3F = 256'h0000FFFFFFFFFFFFFFDF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFF;

DPB dpb_inst_8 (
    .DOA({dpb_inst_8_douta_w[14:0],dpb_inst_8_douta[7]}),
    .DOB({dpb_inst_8_doutb_w[14:0],dpb_inst_8_doutb[7]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({gw_gnd,gw_gnd,ada[14]}),
    .BLKSELB({gw_gnd,gw_gnd,adb[14]}),
    .ADA(ada[13:0]),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[7]}),
    .ADB(adb[13:0]),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[7]})
);

defparam dpb_inst_8.READ_MODE0 = 1'b0;
defparam dpb_inst_8.READ_MODE1 = 1'b1;
defparam dpb_inst_8.WRITE_MODE0 = 2'b00;
defparam dpb_inst_8.WRITE_MODE1 = 2'b00;
defparam dpb_inst_8.BIT_WIDTH_0 = 1;
defparam dpb_inst_8.BIT_WIDTH_1 = 1;
defparam dpb_inst_8.BLK_SEL_0 = 3'b000;
defparam dpb_inst_8.BLK_SEL_1 = 3'b000;
defparam dpb_inst_8.RESET_MODE = "SYNC";
defparam dpb_inst_8.INIT_RAM_00 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_01 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_02 = 256'h0000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_03 = 256'h0000FFFFFFFFFFFFFFFFF415FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_04 = 256'h0000FFFFFFFFFFFFFFFFE595FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_05 = 256'h0000FFFFFFFFFFFFFFFF222EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_06 = 256'h0000FFFFFFFFFFFFFFF9102AF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_07 = 256'h0000FFFFFFFFFFFFFFF411CA5BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_08 = 256'h0000FFFFFFFFFFFFFFFC085C4AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_09 = 256'h0000FFFFFFFFFFFFFFF8C4AC0ABFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0A = 256'h0000FFFFFFFFFFFFFFF94C79D2B7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0B = 256'h0000FFFFFFFFFFFFFFE10572917FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0C = 256'h0000FFFFFFFFFFFFFFE412F401CF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0D = 256'h0000FFFFFFFFFFFFFFC02164A193BFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0E = 256'h0000FFFFFFFFFFFFFFCA21530011FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_0F = 256'h0000FFFFFFFFFFFFFF9AC95412223D2FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_10 = 256'h0000FFFFFFFFFFFFFF1823C0320D3D7BF77F75DBFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_11 = 256'h0000FFFFFFFFFFFFFF11459142507B790485EF6EFFEEDD7C3FFFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_12 = 256'h0000FFFFFFFFFFFFFE20AE5CC4C33670624100040044EFFDD6EFFFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_13 = 256'h0000FFFFFFFFFFFFFC552F18C5203BE01D8048A810510048821FDFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_14 = 256'h0000FFFFFFFFFFFFF883AE2980A266F025C895225A121D9048CADFFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_15 = 256'h0000FFFFFFFFFFFFF8951D312D913C7022219D8213D21A09A8415FFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_16 = 256'h0000FFFFFFFFFFFFF5097D5110265EF0294431A2E146E5D5C1017FFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_17 = 256'h0000FFFFFFFFFFFFE3127C2210D0FCA88126CDDDD526AF22C9814FFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_18 = 256'h0000FFFFFFFFFFFFC522DC862341CA604513326A1CFD847CD20167FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_19 = 256'h0000FFFFFFFFFFFFC82668A20C48DBE01525ADAD5DAA6AB224815FFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_1A = 256'h0000FFFFFFFFFFFFAC02F1844402FDC02385D0E6DA7AFD5675114FFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_1B = 256'h0000FFFFFFFFFFFF3CA4A2248005B5E042C5E45E9EA25BDEB48057FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_1C = 256'h0000FFFFFFFFFFFF38ABF30000A1BDC04A54B4DAD22ADDFD492073FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_1D = 256'h0000FFFFFFFFFFFE4005E1C14182D3D055BF11DBC2ADBE5ED2A123FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_1E = 256'h0000FFFFFFFFFFFC0021D5C0005A62C237DAAD153BB46F57D9D02BFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_1F = 256'h0000FFFFFFFFFFF91215D5953C073E8132A56B5B546C2C595840F3FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_20 = 256'h0000FFFFFFFFFFF9A22B8C82B49763C222532A2225EDBBB4F6B81DFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_21 = 256'h0000FFFFFFFFFFF202D5452120C65683C3ADB25D242BF222DDA039FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_22 = 256'h0000FFFFFFFFFFE30E5D1248C40D67809247CBB6EB9ACD9E65A015FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_23 = 256'h0000FFFFFFFFFFC4847E5C81494FEF02E443ADDA2D558B372AB01EFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_24 = 256'h0000FFFFFFFFFFC452BD225E6C9FCF0A4A6DC5B9B47BAA259A441FFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_25 = 256'h0000FFFFFFFFFF04256D1511929BB7002DE6996A777D9CB3DA41157FFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_26 = 256'h0000FFFFFFFFFF0425585C8819B9BA01115ACCA556D9535A5452197FFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_27 = 256'h0000FFFFFFFFFC2955B24421853DDB011156A41A1D6E262BA8490D7FFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_28 = 256'h0000FFFFFFFFFC204CF24952D8BF5A400A4425277DE902A3D29817BFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_29 = 256'h0000FFFFFFFFFE42AD316D100A3FAFDAD4D100222C1AC444159C0BBFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_2A = 256'h0000FFFFFFFFFEB913619C442176626BFAEFFFEF7FFFA5A000225FFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_2B = 256'h0000FFFFFFFFFEF1FEFA53E50F6B4440100884DF75B7D6ED3A5DA5FFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_2C = 256'h0000FFFFFFFFFF7DFFBE1C694076B4B1228A447779BFD84A01D22F5FFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_2D = 256'h0000FFFFFFFFFFFD7FEFC2A2C0E5F2924C0A8E7FF93BBC92B0284ABFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_2E = 256'h0000FFFFFFFFFFFE7FFDF08481DE5865C626613BE81AD489114522EFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_2F = 256'h0000FFFFFFFFFFFF3FFFDD6221FFF9AB65A5B52DE9177AA480041ADFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_30 = 256'h0000FFFFFFFFFFEFDFFFEB9A05EBDA19EE26533E2C15A64210711357FFFFFFFF;
defparam dpb_inst_8.INIT_RAM_31 = 256'h0000FFFFFFFFFFFFCFFFFFD211DDB86A4621533FE73F4A0C082001F7FFFFFFFF;
defparam dpb_inst_8.INIT_RAM_32 = 256'h0000FFFFFFFFFFFBEFFFFE7A43BDA2BADC12A33ED734BE269C2580DFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_33 = 256'h0000FFFFFFFFFFFDF7FFFFDEA59DF2E0AE05001C47FDC202281081DFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_34 = 256'h0000FFFFFFFFFFFFF9FFFFEFA3BAFBDBCC1DC21E618B5EA29C30AC77FFFFFFFF;
defparam dpb_inst_8.INIT_RAM_35 = 256'h0000FFFFFFFFFFFFF9FFFFFD57BBE44D5C24A23EED9DBB009821A4DBFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_36 = 256'h0000FFFFFFFFFFFFFCFFFFFF7FB6B6925C9BBE37DD99DD094C1920DBFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_37 = 256'h0000FFFFFFFFFFFFDF7FFFFFDF63A2B46E1BA03F64A9D1008C2204BDFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_38 = 256'h0000FFFFFFFFFFFFDF3FFFFFFF6EFA008212D53FB40BFD2A2C1220FDFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_39 = 256'h0000FFFFFFFFFFFFF7DFFFFFFF75FBFFFFFFFFFFFFA3FF204A220A77FFFFFFFF;
defparam dpb_inst_8.INIT_RAM_3A = 256'h0000FFFFFFFFFFFFFFEFFFFFFFFFFFFFE7E6FFFFFFFDFEDFFFBDF3EFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_3B = 256'h0000FFFFFFFFFFFFFFE7FFFF7FFFFFFFFFFFFFFFFFFDFFF91BFF7BDFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_3C = 256'h0000FFFFFFFFFFFFFFF1FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_3D = 256'h0000FFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_3E = 256'h0000FFFFFFFFFFFFFF7EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBFFFFFFFFF;
defparam dpb_inst_8.INIT_RAM_3F = 256'h0000FFFFFFFFFFFFFFFF3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFFFFFFF;

DPB dpb_inst_9 (
    .DOA({dpb_inst_9_douta_w[11:0],dpb_inst_9_douta[7:4]}),
    .DOB({dpb_inst_9_doutb_w[11:0],dpb_inst_9_doutb[7:4]}),
    .CLKA(clka),
    .OCEA(ocea),
    .CEA(cea),
    .RESETA(reseta),
    .WREA(wrea),
    .CLKB(clkb),
    .OCEB(oceb),
    .CEB(ceb),
    .RESETB(resetb),
    .WREB(wreb),
    .BLKSELA({ada[14],ada[13],ada[12]}),
    .BLKSELB({adb[14],adb[13],adb[12]}),
    .ADA({ada[11:0],gw_gnd,gw_gnd}),
    .DIA({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dina[7:4]}),
    .ADB({adb[11:0],gw_gnd,gw_gnd}),
    .DIB({gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,gw_gnd,dinb[7:4]})
);

defparam dpb_inst_9.READ_MODE0 = 1'b0;
defparam dpb_inst_9.READ_MODE1 = 1'b1;
defparam dpb_inst_9.WRITE_MODE0 = 2'b00;
defparam dpb_inst_9.WRITE_MODE1 = 2'b00;
defparam dpb_inst_9.BIT_WIDTH_0 = 4;
defparam dpb_inst_9.BIT_WIDTH_1 = 4;
defparam dpb_inst_9.BLK_SEL_0 = 3'b100;
defparam dpb_inst_9.BLK_SEL_1 = 3'b100;
defparam dpb_inst_9.RESET_MODE = "SYNC";
defparam dpb_inst_9.INIT_RAM_00 = 256'hFFFFFFFFFFFFFFFFEFFFB7DFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_01 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_02 = 256'hFFFFFFFFFFF5FFFFF0DFFFDFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_03 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_04 = 256'hFFFFFFFFFFFFFFFFDFFFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_05 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_06 = 256'hFFFFFFFFFFFFAFFFF70AFFFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_07 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_08 = 256'hFFFFFFFFFFFFFFFFFFEBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_09 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_0A = 256'hFFFFFFFFFFFFF9FFFF70AFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_0B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_0C = 256'hFFFFFFFFFFFFFE7FFD7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_0D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_0E = 256'hFFFFFFFFFFFFFFCFFFFD09FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_0F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_10 = 256'hFFFFFFFFFFFFEFFF5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_11 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_12 = 256'hFFFFFFFFFFFFFFF5FFFF60AFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_13 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_14 = 256'hFFFFFFFFFFBFFBFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_15 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_16 = 256'hFFFFFFFFFFFFFFFFBFFFFB28FFFFFF7FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_17 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_18 = 256'hFFFFFFFFEFFBFFC3FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_19 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_1A = 256'hFFFFFFFFFFFFFFFFF5FFFFF0AFFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_1B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_1C = 256'hFFFFFA53132E82FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_1D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_1E = 256'hFFFFFFFFFFFFFFFFFFDFFFFB2CFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_1F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_20 = 256'hFFFF668181407FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_21 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_22 = 256'hFFFFFFFFFFFFFFFFFFF7EFFF704FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF;
defparam dpb_inst_9.INIT_RAM_23 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_24 = 256'hFFFA25F4D3E0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_25 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7EFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_26 = 256'hFFFFFFFFFFFFFFFFFFFFBEFFFF05FFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_27 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_28 = 256'hFFFFFEFB7DBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_29 = 256'hFFFFFFFFFFFFFFFFFFFEFFFFFFBFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFF;
defparam dpb_inst_9.INIT_RAM_2A = 256'hFFFFFFFFFFFFFFFFFFFFF7DFFFB0EF7DFFFFFFFFFFFFFEFFFFFFFFFFFFBFFFFF;
defparam dpb_inst_9.INIT_RAM_2B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_2C = 256'hFFFFFB7E5FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_2D = 256'hFFDFFFFFFFFF7FFFFFFFFFFFFFFFFFFFFFEFFFFFFFBFFFFFFFFFFF7FFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_2E = 256'hFFFFFFFFFFFFFFFFFFFFFF7DFFF724FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_2F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_30 = 256'hD9B5347FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_31 = 256'hFFFFFFFF7FFFFFFFEFFFFFFFFFFFFFFFFFFFFFFEFEFEFECEEFEEECFDDDBF9F9D;
defparam dpb_inst_9.INIT_RAM_32 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFBFFFF05FFFEFFFFFFFFDFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_33 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_34 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_35 = 256'hFFFFFFFFF7FEFFFDFFFBFFFFFFFFFFFFFBFFFFFFEBFFFFFFFFFDFBFFFFFFFBFF;
defparam dpb_inst_9.INIT_RAM_36 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEFFF09FFFFFFFDFFFFFBFFFFFFFFFDFBFF;
defparam dpb_inst_9.INIT_RAM_37 = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_38 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_39 = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3A = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3B = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3C = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3D = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3E = 256'hFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;
defparam dpb_inst_9.INIT_RAM_3F = 256'h0000000000000000FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF;

DFFE dff_inst_0 (
  .Q(dff_q_0),
  .D(ada[14]),
  .CLK(clka),
  .CE(cea_w)
);
DFFE dff_inst_1 (
  .Q(dff_q_1),
  .D(adb[14]),
  .CLK(clkb),
  .CE(ceb_w)
);
DFFE dff_inst_2 (
  .Q(dff_q_2),
  .D(dff_q_1),
  .CLK(clkb),
  .CE(oceb)
);
MUX2 mux_inst_4 (
  .O(douta[0]),
  .I0(dpb_inst_0_douta[0]),
  .I1(dpb_inst_4_douta[0]),
  .S0(dff_q_0)
);
MUX2 mux_inst_9 (
  .O(douta[1]),
  .I0(dpb_inst_1_douta[1]),
  .I1(dpb_inst_4_douta[1]),
  .S0(dff_q_0)
);
MUX2 mux_inst_14 (
  .O(douta[2]),
  .I0(dpb_inst_2_douta[2]),
  .I1(dpb_inst_4_douta[2]),
  .S0(dff_q_0)
);
MUX2 mux_inst_19 (
  .O(douta[3]),
  .I0(dpb_inst_3_douta[3]),
  .I1(dpb_inst_4_douta[3]),
  .S0(dff_q_0)
);
MUX2 mux_inst_24 (
  .O(douta[4]),
  .I0(dpb_inst_5_douta[4]),
  .I1(dpb_inst_9_douta[4]),
  .S0(dff_q_0)
);
MUX2 mux_inst_29 (
  .O(douta[5]),
  .I0(dpb_inst_6_douta[5]),
  .I1(dpb_inst_9_douta[5]),
  .S0(dff_q_0)
);
MUX2 mux_inst_34 (
  .O(douta[6]),
  .I0(dpb_inst_7_douta[6]),
  .I1(dpb_inst_9_douta[6]),
  .S0(dff_q_0)
);
MUX2 mux_inst_39 (
  .O(douta[7]),
  .I0(dpb_inst_8_douta[7]),
  .I1(dpb_inst_9_douta[7]),
  .S0(dff_q_0)
);
MUX2 mux_inst_44 (
  .O(doutb[0]),
  .I0(dpb_inst_0_doutb[0]),
  .I1(dpb_inst_4_doutb[0]),
  .S0(dff_q_2)
);
MUX2 mux_inst_49 (
  .O(doutb[1]),
  .I0(dpb_inst_1_doutb[1]),
  .I1(dpb_inst_4_doutb[1]),
  .S0(dff_q_2)
);
MUX2 mux_inst_54 (
  .O(doutb[2]),
  .I0(dpb_inst_2_doutb[2]),
  .I1(dpb_inst_4_doutb[2]),
  .S0(dff_q_2)
);
MUX2 mux_inst_59 (
  .O(doutb[3]),
  .I0(dpb_inst_3_doutb[3]),
  .I1(dpb_inst_4_doutb[3]),
  .S0(dff_q_2)
);
MUX2 mux_inst_64 (
  .O(doutb[4]),
  .I0(dpb_inst_5_doutb[4]),
  .I1(dpb_inst_9_doutb[4]),
  .S0(dff_q_2)
);
MUX2 mux_inst_69 (
  .O(doutb[5]),
  .I0(dpb_inst_6_doutb[5]),
  .I1(dpb_inst_9_doutb[5]),
  .S0(dff_q_2)
);
MUX2 mux_inst_74 (
  .O(doutb[6]),
  .I0(dpb_inst_7_doutb[6]),
  .I1(dpb_inst_9_doutb[6]),
  .S0(dff_q_2)
);
MUX2 mux_inst_79 (
  .O(doutb[7]),
  .I0(dpb_inst_8_doutb[7]),
  .I1(dpb_inst_9_doutb[7]),
  .S0(dff_q_2)
);
endmodule //blk_mem_gen_4
